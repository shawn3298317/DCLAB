//*************************************************************************************************//
// File: exp1_traffic.v                                                                            //
// Description: This is the verilog file for traffic light control logic                           //
//*************************************************************************************************//



//*  
// @parameter clk   : 50MHz clock signal
// @parameter reset : reset signal
// @parameter change: change signal
//*
module traffic_ctr (
	clk,
	reset,
	change
	);
	

//*******combinational part*********//





//*******sequential part************//

	
	
endmodule

